module ALUControl(ALUOp, instr5_0, ALUCntrl);
  
